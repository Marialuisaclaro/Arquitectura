library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address   : in  std_logic_vector(11 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (

"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000000", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000001", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000011", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000010", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000011", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000011", --('MOV', '(Dir)', 'A')
"000010110100000000000000001100000011", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000100", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000101", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000110", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000111", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000001000", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000001001", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000001010", --('MOV', '(Dir)', 'A')
"000010110100000000000101010101010101", --('MOV', 'A', 'Lit')
"000000001100000101000000000000001011", --('MOV', '(Dir)', 'A')
"000010110100000000001010101010101010", --('MOV', 'A', 'Lit')
"000000001100000101000000000000001100", --('MOV', '(Dir)', 'A')
"000100000000010011010000000001111010", --('CALL', 'INS')
"000100000000010011010000000001111010", --('CALL', 'INS')
"000001110100000000000000000000001000", --('MOV', 'B', 'Lit')
"000000101100001101000000000000000000", --('IN', '(B)', 'Lit')
"000100000000010011010000000001111010", --('CALL', 'INS')
"000001110100000000000000000000001001", --('MOV', 'B', 'Lit')
"000000101100001101000000000000000000", --('IN', '(B)', 'Lit')
"000010111000000000000000000000000100", --('MOV', 'A', '(Dir)')
"001000000100000000000000000000000000", --('OUT', 'A', 'Lit')
"000100000000010011010000000000101100", --('CALL', 'INS')
"000010111000000000000000000000000011", --('MOV', 'A', '(Dir)')
"000000000100100000000000000000000000", --('CMP', 'A', 'Lit')
"001100000000000010000000000001011110", --('JEQ', 'INS')
"000100000000010011010000000001000100", --('CALL', 'INS')
"000010111000000000000000000000000010", --('MOV', 'A', '(Dir)')
"000000000100100000000000000000000000", --('CMP', 'A', 'Lit')
"001100000000000010000000000001011110", --('JEQ', 'INS')
"000100000000000010000000000000100011", --('JMP', 'INS')
"000010111000000000000000000000000110", --('MOV', 'A', '(Dir)')
"001000000100000000000000000000000001", --('OUT', 'A', 'Lit')
"000100000000010011010000000001111010", --('CALL', 'INS')
"000001110100000000000000000000000101", --('MOV', 'B', 'Lit')
"000000101100001101000000000000000000", --('IN', '(B)', 'Lit')
"000010111000000000000000000000000110", --('MOV', 'A', '(Dir)')
"000010001001100000000000000000000101", --('OR', 'A', '(Dir)')
"000000001100000101000000000000000110", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000001001", --('MOV', 'A', '(Dir)')
"000010001001000000000000000000000101", --('AND', 'A', '(Dir)')
"000000000100100000000000000000000000", --('CMP', 'A', 'Lit')
"001100000000000010000000000001011100", --('JEQ', 'INS')
"000001001100000000000000000000000000", --('MOV', 'B', 'A')
"000010111000000000000000000000001001", --('MOV', 'A', '(Dir)')
"000010000000100000000000000000000000", --('SUB', 'A', 'B')
"000000001100000101000000000000001001", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000000011", --('MOV', 'A', '(Dir)')
"000010000100100000000000000000000001", --('SUB', 'A', 'Lit')
"000000001100000101000000000000000011", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000000100", --('MOV', 'A', '(Dir)')
"000010000100100000000000000000000001", --('SUB', 'A', 'Lit')
"000000001100000101000000000000000100", --('MOV', '(Dir)', 'A')
"001000000100000000000000000000000000", --('OUT', 'A', 'Lit')
"000100000000000010000000000001011100", --('JMP', 'INS')
"000010111000000000000000000000000111", --('MOV', 'A', '(Dir)')
"001000000100000000000000000000000001", --('OUT', 'A', 'Lit')
"000100000000010011010000000001111010", --('CALL', 'INS')
"000001110100000000000000000000000101", --('MOV', 'B', 'Lit')
"000000101100001101000000000000000000", --('IN', '(B)', 'Lit')
"000010111000000000000000000000000111", --('MOV', 'A', '(Dir)')
"000010001001100000000000000000000101", --('OR', 'A', '(Dir)')
"000000001100000101000000000000000111", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000001000", --('MOV', 'A', '(Dir)')
"000010001001000000000000000000000101", --('AND', 'A', '(Dir)')
"000000000100100000000000000000000000", --('CMP', 'A', 'Lit')
"001100000000000010000000000001011100", --('JEQ', 'INS')
"000001001100000000000000000000000000", --('MOV', 'B', 'A')
"000010111000000000000000000000001000", --('MOV', 'A', '(Dir)')
"000010000000100000000000000000000000", --('SUB', 'A', 'B')
"000000001100000101000000000000001000", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000000010", --('MOV', 'A', '(Dir)')
"000010000100100000000000000000000001", --('SUB', 'A', 'Lit')
"000000001100000101000000000000000010", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000000100", --('MOV', 'A', '(Dir)')
"000010000100100000000000000100000000", --('SUB', 'A', 'Lit')
"000000001100000101000000000000000100", --('MOV', '(Dir)', 'A')
"001000000100000000000000000000000000", --('OUT', 'A', 'Lit')
"000100000000000010000000000001011100", --('JMP', 'INS')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000010110100000000000000001011101110", --('MOV', 'A', 'Lit')
"000100000000010011010000000001100010", --('CALL', 'INS')
"000100000000010011010000000001101110", --('CALL', 'INS')
"000100000000000010000000000001011110", --('JMP', 'INS')
"000000001100010101010000000000000000", --('PUSH', 'A')
"000010000011100000000000000000000000", --('SHR', 'A')
"000000001100010101010000000000000000", --('PUSH', 'A')
"000010111000000000000000000000001011", --('MOV', 'A', '(Dir)')
"001000000100000000000000000000000001", --('OUT', 'A', 'Lit')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000100000000010011010000000010100111", --('CALL', 'INS')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000001100010101010000000000000000", --('PUSH', 'A')
"000010000011100000000000000000000000", --('SHR', 'A')
"000000001100010101010000000000000000", --('PUSH', 'A')
"000010111000000000000000000000001100", --('MOV', 'A', '(Dir)')
"001000000100000000000000000000000001", --('OUT', 'A', 'Lit')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000100000000010011010000000010100111", --('CALL', 'INS')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000110000010101010000000000000000", --('PUSH', 'B')
"000010101100000000000000000000000001", --('IN', 'A', 'Lit')
"000001101100000000000000000000000001", --('IN', 'B', 'Lit')
"000000000000100000000000000000000000", --('CMP', 'A', 'B')
"001100000000000010000000000001111100", --('JEQ', 'INS')
"000001000010100000000000000000000000", --('XOR', 'B', 'A')
"000010101100000000000000000000000001", --('IN', 'A', 'Lit')
"000010000001000000000000000000000000", --('AND', 'A', 'B')
"000000000100100000000000000000000000", --('CMP', 'A', 'Lit')
"010100000000000010000000000010000000", --('JNE', 'INS')
"000010110000000000000000000000000000", --('MOV', 'A', 'B')
"000000000000000000100000000000000000", --('POP', 'B')
"000001111000010100000000000000000000", --('POP', 'B')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000110000010101010000000000000000", --('PUSH', 'B')
"000001101100000000000000000000000010", --('IN', 'B', 'Lit')
"000000000000100000000000000000000000", --('CMP', 'A', 'B')
"011100000000000010000000000010001010", --('JGT', 'INS')
"000000000000000000100000000000000000", --('POP', 'B')
"000001111000010100000000000000000000", --('POP', 'B')
"000100000000000010000000000010010011", --('JMP', 'INS')
"000001001100000000000000000000000000", --('MOV', 'B', 'A')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000000110000010101010000000000000000", --('PUSH', 'B')
"000001101100000000000000000000000010", --('IN', 'B', 'Lit')
"000000000000100000000000000000000000", --('CMP', 'A', 'B')
"010100000000000010000000000010100011", --('JNE', 'INS')
"000000000000000000100000000000000000", --('POP', 'B')
"000001111000010100000000000000000000", --('POP', 'B')
"000000001100010101010000000000000000", --('PUSH', 'A')
"000010110000000000000000000000000000", --('MOV', 'A', 'B')
"000001101100000000000000000000000011", --('IN', 'B', 'Lit')
"000000000000100000000000000000000000", --('CMP', 'A', 'B')
"011100000000000010000000000010010000", --('JGT', 'INS')
"000001001100000000000000000000000000", --('MOV', 'B', 'A')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000000000000000100000000000000000", --('POP', 'B')
"000001111000010100000000000000000000", --('POP', 'B')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000001100010101010000000000000000", --('PUSH', 'A')
"000000110000010101010000000000000000", --('PUSH', 'B')
"000001101100000000000000000000000011", --('IN', 'B', 'Lit')
"000010000000000000000000000000000000", --('ADD', 'A', 'B')
"000001101100000000000000000000000010", --('IN', 'B', 'Lit')
"000000000100100000000000001111101000", --('CMP', 'A', 'Lit')
"100100000000000010000000000010110001", --('JLT', 'INS')
"000010000100100000000000001111101000", --('SUB', 'A', 'Lit')
"000001010000000000000000000000000001", --('INC', 'B')
"000100000000000010000000000010101100", --('JMP', 'INS')
"000010000010100000000000000000000000", --('XOR', 'A', 'B')
"000001000010100000000000000000000000", --('XOR', 'B', 'A')
"000010000010100000000000000000000000", --('XOR', 'A', 'B')
"000100000000010011010000000010001001", --('CALL', 'INS')
"000000000000000000100000000000000000", --('POP', 'B')
"000001111000010100000000000000000000", --('POP', 'B')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000" --blank
); 
begin
   dataout <= memory(to_integer(unsigned(address))); 
end Behavioral; 

