library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address   : in  std_logic_vector(11 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (
    "000010110100000000000000000000000011",-- MOV A,3
    "000000001100000101000000000000000000",-- MOV (var1),A
    "000010110100000000000000000000000100",-- MOV A,4
    "000000001100000101000000000000000001",-- MOV (var2),A
    "000010110100000000000000000000000000",-- MOV A,0
    "000000001100000101000000000000000010",-- MOV (res),A
    "000010110100000000000000000000000000",-- MOV A,0
    "000000001100000101000000000000000011",-- MOV (i),A
    "000010111000000000000000000000000000",-- MOV A,(var1)     <= start
    "000001111000000000000000000000000011",-- MOV B,(i)
    "000000000000100000000000000000000000",-- CMP A, B
    "001100000000000010000000000000010011", --JEQ save
    "000010111000000000000000000000000010", --MOV A,(res)
    "000010001000000000000000000000000001", --ADD A,(var2)
    "000000001100000101000000000000000010", --MOV (res),A
    "000010111000000000000000000000000011", --MOV A,(i)
    "000010000100000000000000000000000001", --ADD A,1
    "000000001100000101000000000000000011", --MOV (i),A
    "000100000000000010000000000000001000", --JMP start
    "000001111000000000000000000000000010", --MOV B,(res)   <= save
    "000100000000000010000000000000010100", --JMP end       <= end
    "000000000000000000000000000000000000", --39
    "000000000000000000000000000000000000", -- BLANKS
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000", 	 
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000"
        ); 
begin

   dataout <= memory(to_integer(unsigned(address))); 

end Behavioral; 
