library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address   : in  std_logic_vector(11 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (

"000010110100000000000000000000000101", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000000", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000001010", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000001", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000001", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000010", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000011", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000011", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000001000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000100", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000101", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000101", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000110", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000110", --('MOV', '(Dir)', 'A')
"000010110100000000000000000000000000", --('MOV', 'A', 'Lit')
"000000001100000101000000000000000111", --('MOV', '(Dir)', 'A')
"000001110100000000000000000000000000", --('MOV', 'B', 'Lit')
"000010111000000000000000000000000110", --('MOV', 'A', '(Dir)')
"000000000100100000000000000000000000", --('CMP', 'A', 'Lit')
"001100000000000010000000000000100010", --('JEQ', 'INS')
"000010000100100000000000000000000001", --('DEC', 'A')
"000000001100000101000000000000000110", --('MOV', '(Dir)', 'A')
"000010111000000000000000000000000111", --('MOV', 'A', '(Dir)')
"000010001000001000000000000000000000", --('ADD', 'A', '(B)')
"000000001100000101000000000000000111", --('MOV', '(Dir)', 'A')
"000001010000000000000000000000000001", --('INC', 'B')
"000100000000000010000000000000010111", --('JMP', 'INS')
"000010111000000000000000000000000111", --('MOV', 'A', '(Dir)')
"000100000000000010000000000000100010", --('JMP', 'INS')
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000" --blank
); 
begin
   dataout <= memory(to_integer(unsigned(address))); 
end Behavioral; 

