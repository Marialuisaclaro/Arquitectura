library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        address   : in  std_logic_vector(11 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (

"000010110100000000000000000000001011", --('MOV', 'A', 'Lit')
"000001110100000000000000000000010101", --('MOV', 'B', 'Lit')
"000000001100010101010000000000000000", --('PUSH', 'A')
"000000110000010101010000000000000000", --('PUSH', 'B')
"000000000000000000100000000000000000", --('POP', 'A')
"000010111000010100000000000000000000", --('POP', 'A')
"000000000000000000100000000000000000", --('POP', 'B')
"000001111000010100000000000000000000", --('POP', 'B')
"000100000000010011010000000000001011", --('CALL', 'INS')
"000001000000000000000000000000000000", --('ADD', 'B', 'A')
"000100000000000010000000000000001010", --('JMP', 'INS')
"000010000000000000000000000000000000", --('ADD', 'A', 'B')
"000000000000000000100000000000000000", --RET
"000100000000010000000000000000000000", --RET
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000", --blank
"000000000000000000000000000000000000" --blank
); 
begin
   dataout <= memory(to_integer(unsigned(address))); 
end Behavioral; 

